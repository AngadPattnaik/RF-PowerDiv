*Including the 180nm technology file
.include 180nm_bulk.txt
.option rshunt = 1.0e12

vgg1 6 3 dc 1.4v
m1 1 6 3 0 NMOS W=80u
vdd1 1 10 dc 0.6v
ld1 10 3 100n

vgg2 4 b dc 1.4v
m2 c 4 b 0 NMOS W=80u 
vdd2 c 11 dc 0.6v
ld2 11 b 100n

vgg3 5 2 dc 1.4v
m3 a 5 2 0 NMOS W=80u 
vdd3 a 12 dc 0.6v
ld3 12 2 100n

c1 1 9 1n
c2 a 7 1n
c3 b 8 1n

csa 3 a 1n
csb 2 b 1n
csc 1 c 1n

V1 10 0 dc 0 ac 1 

r1 9 10 50
r2 7 0 50
r3 8 0 50
.ac dec 10  100Meg 100G

.control
run

plot vdb(7) vdb(8) xlog

*plot {57.29*vp(7)} {57.29*vp(8)} xlog

.endc

.end



