*Including the 180nm technology file
.include 180nm_bulk.txt
.option rshunt = 1.0e12


m1 1 6 3 0 NMOS W=80u m=12
vgg1 p 0 dc 1.4v
la 6 p 100n
vdd1 10 0 dc 0.8v
ld1 1 10 100n

m2 c 4 b 0 NMOS W=80u m=12 
vgg2 l 0 dc 1.4v
lb 4 l 100n
vdd2 11 0 dc 0.8v
ld2 c 11 100n

m3 a 5 2 0 NMOS W=80u m=12 
vgg3 m 0 dc 1.4v
lc 5 m 100n
vdd3 12 0 dc 0.8v
ld3 a 12 100n


c2 a 7 10n
c3 b 8 10n
r2 7 0 50
r3 8 0 50

csa 3 a 10n
csb 2 b 10n
csc 1 c 10n


c1 1 9 10n

V1 9 0 dc 0 ac 1 


.ac dec 10  100Meg 500G

.control
run

plot vdb(7) vdb(8) xlog
print vdb(7)



.endc

.end



